library verilog;
use verilog.vl_types.all;
entity fabrica_vlg_vec_tst is
end fabrica_vlg_vec_tst;
