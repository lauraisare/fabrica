library verilog;
use verilog.vl_types.all;
entity fabrica_vlg_check_tst is
    port(
        c               : in     vl_logic;
        d               : in     vl_logic;
        e               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fabrica_vlg_check_tst;
